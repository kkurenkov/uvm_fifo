// ----------------------------------------------------------------------------
// Author:   Konstantin Kurenkov
// Email:    krendkrend@gmail.com
// FileName: kvt_scfifo_tb_inc.sv
// Create date: 16/11/2021
//
// Description: Main Include files for SCFIFO Example
//
// ----------------------------------------------------------------------------

`include "uvm_macros.svh"
`include "kvt_scfifo_env_pkg.sv"

import uvm_pkg::*;
import kvt_scfifo_env_pkg::*;

`include "kvt_scfifo_wrapper.sv"
`include "kvt_scfifo_tb_top.sv"